entity ( 
    port(
        --comentario
        --x2
        --x3
    )
)