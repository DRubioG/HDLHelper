entity hola is
end entity hola;

